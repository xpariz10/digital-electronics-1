library ieee;
use ieee.std_logic_1164.all;

entity s_debouncing is
  Generic(
    clk_f	    : integer := 50_000_000;  --system clock frequency in Hz
    wait_time : integer := 120);        --time to wait in ms
  Port(
    clk     : in  std_logic;  
    rst	    : in  std_logic;  
    button  : in  std_logic;
    en      : in  std_logic;
    result  : out std_logic); 
end s_debouncing;

architecture Behavioral of s_debouncing is
begin
    
clk_enable : entity work.clk_en_db
      port map (
          clk => clk,
          rst => rst,
          ce   => en
      );
    
    p_s_debouncing : process (clk, rst) is
    begin
        if rising_edge(clk) then
           	if (rst = '1') then
               	result <= '0';
           	elsif (button = '1' and en = '1')
           		result <= '1';
            else
            	result <= '0';
       		end if;
        end if;
    end process p_d_ff_rst;
end architecture Behavioral;
